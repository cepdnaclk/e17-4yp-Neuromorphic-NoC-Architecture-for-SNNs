`timescale 1ns/100ps

module pr_id_ex (
    CLK, RESET, 

    ID_PC, ID_REG_DATA1, ID_REG_DATA2, ID_IMMEDIATE,
    ID_REG_WRITE_ADDR, ID_REG_READ_ADDR1, ID_REG_READ_ADDR2, 
    ID_ALU_SELECT, ID_OPERAND1_SELECT, ID_OPERAND2_SELECT,
    ID_REG_WRITE_EN, ID_DATA_MEM_WRITE, ID_DATA_MEM_READ, 
    ID_BRANCH_CTRL, ID_WB_VALUE_SELECT,

    EX_PC, EX_REG_DATA1, EX_REG_DATA2, EX_IMMEDIATE,
    EX_REG_WRITE_ADDR, EX_REG_READ_ADDR1, EX_REG_READ_ADDR2,
    EX_ALU_SELECT, EX_OPERAND1_SELECT, EX_OPERAND2_SELECT,
    EX_REG_WRITE_EN, EX_DATA_MEM_WRITE, EX_DATA_MEM_READ,
    EX_BRANCH_CTRL, EX_WB_VALUE_SELECT
);

    input CLK, RESET;

    input [31:0] ID_PC, ID_REG_DATA1, ID_REG_DATA2, ID_IMMEDIATE;
    input [4:0] ID_REG_WRITE_ADDR, ID_REG_READ_ADDR1, ID_REG_READ_ADDR2;
    input ID_REG_WRITE_EN, ID_OPERAND1_SELECT, ID_OPERAND2_SELECT;
    input [5:0] ID_ALU_SELECT;
    input [3:0] ID_DATA_MEM_READ, ID_BRANCH_CTRL;
    input [2:0] ID_DATA_MEM_WRITE;
    input [1:0] ID_WB_VALUE_SELECT;

    output reg [31:0] EX_PC, EX_REG_DATA1, EX_REG_DATA2, EX_IMMEDIATE;
    output reg [4:0] EX_REG_WRITE_ADDR, EX_REG_READ_ADDR1, EX_REG_READ_ADDR2;
    output reg EX_REG_WRITE_EN, EX_OPERAND1_SELECT, EX_OPERAND2_SELECT;
    output reg [5:0] EX_ALU_SELECT;
    output reg [3:0] EX_DATA_MEM_READ, EX_BRANCH_CTRL;
    output reg [2:0] EX_DATA_MEM_WRITE;
    output reg [1:0] EX_WB_VALUE_SELECT;

    always @ (posedge CLK)
    begin
        #1
        if (RESET == 1'b1)
        begin
            EX_PC = 32'b0;
            EX_REG_DATA1 = 32'b0;
            EX_REG_DATA2 = 32'b0;
            EX_IMMEDIATE = 32'b0;
            EX_REG_WRITE_ADDR = 4'b0;
            EX_REG_READ_ADDR1 = 4'b0;
            EX_REG_READ_ADDR2 = 4'b0;
            EX_ALU_SELECT = 5'b0;
            EX_OPERAND1_SELECT = 1'b0;
            EX_OPERAND2_SELECT = 1'b0;
            EX_REG_WRITE_EN = 1'b0;
            EX_DATA_MEM_WRITE = 3'b0;
            EX_DATA_MEM_READ = 4'b0;
            EX_BRANCH_CTRL = 4'b0;
            EX_WB_VALUE_SELECT = 2'b0;
        end
        else
        begin
            EX_PC = ID_PC;
            EX_REG_DATA1 = ID_REG_DATA1;
            EX_REG_DATA2 = ID_REG_DATA2;
            EX_IMMEDIATE = ID_IMMEDIATE;
            EX_REG_WRITE_ADDR = ID_REG_WRITE_ADDR;
            EX_REG_READ_ADDR1 = ID_REG_READ_ADDR1;
            EX_REG_READ_ADDR2 = ID_REG_READ_ADDR2;
            EX_ALU_SELECT = ID_ALU_SELECT;
            EX_OPERAND1_SELECT = ID_OPERAND1_SELECT;
            EX_OPERAND2_SELECT = ID_OPERAND2_SELECT;
            EX_REG_WRITE_EN = ID_REG_WRITE_EN;
            EX_DATA_MEM_WRITE = ID_DATA_MEM_WRITE;
            EX_DATA_MEM_READ = ID_DATA_MEM_READ;
            EX_BRANCH_CTRL = ID_BRANCH_CTRL;
            EX_WB_VALUE_SELECT = ID_WB_VALUE_SELECT;
        end
    end
    
endmodule